configuration cfg of SADg_tb is
	for sadg_test
		-- use default configuration
	end for;
end cfg;