configuration cfg of SAD_tb is
	for sad_test
		-- use default configuration
	end for;
end cfg;